covergroup CovKind;

    CP1: coverpoint tr.i
    {
        ignore_bins even = {6,7};
    }

endgroup

/*

*/