/*
    purpose: This file contains example of score board
    Author: Karim Mahmoud Kamal
    Date:    7th of February 2024
*/

module score_board();

    initial begin
        

    end
endmodule

