/*
    purpose: This file contains some tasks examples
    Author: Karim Mahmoud Kamal
    Date:    11th of February 2024
*/

module Function1();

    // Task
    function my_log ( );
        $display("Hello from my_log task");
        $display("Hello from my_log task");
    endfunction

    initial begin
        my_log();
    end

endmodule
