/*
    purpose: This file contains exapmle of top module of adder
    Author: Karim Mahmoud Kamal
    Date:    17th of February 2024
*/

module adder ( intf.dut abc );
    assign abc.c = abc.a + abc.b;
endmodule