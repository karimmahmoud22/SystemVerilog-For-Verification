/*
    purpose: This file contains exapmle of interface
    Author: Karim Mahmoud Kamal
    Date:    17th of February 2024
*/

interface arb_int( input bit clk );
    logic [1:0] request, grant;
    logic rst;

endinterface
