/*
    purpose: This file contains example of ATM Router header with interface
    Author: Karim Mahmoud Kamal
    Date:    23th of February 2024
*/

module atm_router(
    Rx_if.DUT Rx0, Rx1, Rx2, Rx3,
    Tx_if.DUT Tx0, Tx1, Tx2, Tx3,
    input logic clk, rst);

endmodule