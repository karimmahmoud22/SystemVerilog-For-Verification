/*
    purpose: This file contains how to disable implicit nets in SystemVerilog
    Author: Karim Mahmoud Kamal
    Date:    15th of February 2024
*/

// To disable implicit nets in SystemVerilog, use the following line
'default_nettype none

module casting();

endmodule

