/*
    purpose: This file contains example of environment using mailbox
    Author: Karim Mahmoud Kamal
    Date:    25th of April 2024
*/