module designx (intf.dut abc);
    initial begin
        abc.addr <= 8'hFF;
    end
endmodule