covergroup SequenceOfTransitions;
    coverpoint a {
        bins t1 = ( 0 => 1 ) , ( 0 => 2) , ( 0 => 3);
    }
    
endgroup