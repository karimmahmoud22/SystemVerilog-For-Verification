covergroup CovKind;

    kind: coverpoint tr.kind;
    port: coverpoint tr.port;
    cross kind, port;

endgroup

/*

*/