bit running =1;

module bus ( bus_interface.dut abc );

endmodule